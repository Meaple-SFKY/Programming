module aluMod (
	input wire clk,
	input wire [5:0] funct,
	input wire [31:0] muxSecOut, muxThiOut,
	output reg [31:0] aluOut
);
	
	always @(posedge clk) begin
		
	end

endmodule