module ctrlUniMod (
	input wire clk, rst,
	input wire [5:0] irOutOpe,
	output wire ifWR, wriReg, muxSegSig, muxThiSig, funct, datMemWr, wbSig
);
	
endmodule